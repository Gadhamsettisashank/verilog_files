module tb_decoder2to4;

    reg [1:0] in;
    reg en;
    wire [3:0] out;

    decoder2to4 uut (
        .in(in),
        .en(en),
        .out(out)
    );

    initial begin
        $display("Time | en in | out");
        $monitor("%4t | %b  %b  | %b", $time, en, in, out);

        en = 0; in = 2'b00; #10;
        en = 1; in = 2'b00; #10;
        in = 2'b01; #10;
        in = 2'b10; #10;
        in = 2'b11; #10;
        en = 0; #10;

        $finish;
    end

endmodule
